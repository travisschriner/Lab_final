----------------------------------------------------------------------------------
-- Company: USAFA DFEC
-- Engineer: C2C Travis Schriner
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity LUT is
	port( val 	: in unsigned (7 downto 0);
			level : out unsigned(7 downto 0)
		 );
end LUT;

architecture Behavioral of LUT is

begin
process(val)
begin
	case val is
		when ("00000000") =>
			level <= ("00000000");
		when to_unsigned(1, 8) =>
			level <= to_unsigned(2, 8);
		when to_unsigned(2, 8) =>
			level <= to_unsigned(4, 8);
		when to_unsigned(3, 8) =>
			level <= to_unsigned(6, 8);
		when to_unsigned(4, 8) =>
			level <= to_unsigned(8, 8);
		when to_unsigned(5, 8) =>
			level <= to_unsigned(10, 8);
		when to_unsigned(6, 8) =>
			level <= to_unsigned(12, 8);
		when to_unsigned(7, 8) =>
			level <= to_unsigned(14, 8);
		when to_unsigned(8, 8) =>
			level <= to_unsigned(16, 8);
		when to_unsigned(9, 8) =>
			level <= to_unsigned(18, 8);
		when to_unsigned(10, 8) =>
			level <= to_unsigned(20, 8);
		when to_unsigned(11, 8) =>
			level <= to_unsigned(22, 8);
		when to_unsigned(12, 8) =>
			level <= to_unsigned(24, 8);
		when to_unsigned(13, 8) =>
			level <= to_unsigned(26, 8);
		when to_unsigned(14, 8) =>
			level <= to_unsigned(28, 8);
		when to_unsigned(15, 8) =>
			level <= to_unsigned(30, 8);
		when to_unsigned(16, 8) =>
			level <= to_unsigned(32, 8);
		when to_unsigned(17, 8) =>
			level <= to_unsigned(34, 8);
		when to_unsigned(18, 8) =>
			level <= to_unsigned(36, 8);
		when to_unsigned(19, 8) =>
			level <= to_unsigned(38, 8);
		when to_unsigned(20, 8) =>
			level <= to_unsigned(40, 8);
		when to_unsigned(21, 8) =>
			level <= to_unsigned(42, 8);
		when to_unsigned(22, 8) =>
			level <= to_unsigned(44, 8);
		when to_unsigned(23, 8) =>
			level <= to_unsigned(46, 8);
		when to_unsigned(24, 8) =>
			level <= to_unsigned(48, 8);
		when to_unsigned(25, 8) =>
			level <= to_unsigned(50, 8);
		when to_unsigned(26, 8) =>
			level <= to_unsigned(52, 8);
		when to_unsigned(27, 8) =>
			level <= to_unsigned(54, 8);
		when to_unsigned(28, 8) =>
			level <= to_unsigned(56, 8);
		when to_unsigned(29, 8) =>
			level <= to_unsigned(58, 8);
		when to_unsigned(30, 8) =>
			level <= to_unsigned(60, 8);
		when to_unsigned(31, 8) =>
			level <= to_unsigned(62, 8);
		when to_unsigned(32, 8) =>
			level <= to_unsigned(66, 8);
		when to_unsigned(33, 8) =>
			level <= to_unsigned(68, 8);
		when to_unsigned(34, 8) =>
			level <= to_unsigned(70, 8);
		when to_unsigned(35, 8) =>
			level <= to_unsigned(72, 8);
		when to_unsigned(36, 8) =>
			level <= to_unsigned(74, 8);
		when to_unsigned(37, 8) =>
			level <= to_unsigned(76, 8);
		when to_unsigned(38, 8) =>
			level <= to_unsigned(78, 8);
		when to_unsigned(39, 8) =>
			level <= to_unsigned(80, 8);
		when to_unsigned(40, 8) =>
			level <= to_unsigned(82, 8);
		when to_unsigned(41, 8) =>
			level <= to_unsigned(84, 8);
		when to_unsigned(42, 8) =>
			level <= to_unsigned(86, 8);
		when to_unsigned(43, 8) =>
			level <= to_unsigned(88, 8);
		when to_unsigned(44, 8) =>
			level <= to_unsigned(90, 8);
		when to_unsigned(45, 8) =>
			level <= to_unsigned(92, 8);
		when to_unsigned(46, 8) =>
			level <= to_unsigned(94, 8);
		when to_unsigned(47, 8) =>
			level <= to_unsigned(96, 8);
		when to_unsigned(48, 8) =>
			level <= to_unsigned(98, 8);
		when to_unsigned(49, 8) =>
			level <= to_unsigned(100, 8);
		when to_unsigned(50, 8) =>
			level <= to_unsigned(102, 8);
		when to_unsigned(51, 8) =>
			level <= to_unsigned(104, 8);
		when to_unsigned(52, 8) =>
			level <= to_unsigned(106, 8);
		when to_unsigned(53, 8) =>
			level <= to_unsigned(108, 8);
		when to_unsigned(54, 8) =>
			level <= to_unsigned(110, 8);
		when to_unsigned(55, 8) =>
			level <= to_unsigned(112, 8);
		when to_unsigned(56, 8) =>
			level <= to_unsigned(114, 8);
		when to_unsigned(57, 8) =>
			level <= to_unsigned(116, 8);
		when to_unsigned(58, 8) =>
			level <= to_unsigned(118, 8);
		when to_unsigned(59, 8) =>
			level <= to_unsigned(120, 8);
		when to_unsigned(60, 8) =>
			level <= to_unsigned(122, 8);
		when to_unsigned(61, 8) =>
			level <= to_unsigned(124, 8);
		when to_unsigned(62, 8) =>
			level <= to_unsigned(126, 8);
		when to_unsigned(63, 8) =>
			level <= to_unsigned(128, 8);
		when to_unsigned(64, 8) =>
			level <= to_unsigned(130, 8);
		when to_unsigned(65, 8) =>
			level <= to_unsigned(132, 8);
		when to_unsigned(66, 8) =>
			level <= to_unsigned(134, 8);
		when to_unsigned(67, 8) =>
			level <= to_unsigned(136, 8);
		when to_unsigned(68, 8) =>
			level <= to_unsigned(138, 8);
		when to_unsigned(69, 8) =>
			level <= to_unsigned(140, 8);
		when to_unsigned(70, 8) =>
			level <= to_unsigned(142, 8);
		when to_unsigned(71, 8) =>
			level <= to_unsigned(144, 8);
		when to_unsigned(72, 8) =>
			level <= to_unsigned(146, 8);
		when to_unsigned(73, 8) =>
			level <= to_unsigned(148, 8);
		when to_unsigned(74, 8) =>
			level <= to_unsigned(150, 8);
		when to_unsigned(75, 8) =>
			level <= to_unsigned(152, 8);
		when to_unsigned(76, 8) =>
			level <= to_unsigned(154, 8);
		when to_unsigned(77, 8) =>
			level <= to_unsigned(156, 8);
		when to_unsigned(78, 8) =>
			level <= to_unsigned(158, 8);
		when to_unsigned(79, 8) =>
			level <= to_unsigned(160, 8);
		when to_unsigned(80, 8) =>
			level <= to_unsigned(162, 8);
		when to_unsigned(81, 8) =>
			level <= to_unsigned(164, 8);
		when to_unsigned(82, 8) =>
			level <= to_unsigned(166, 8);
		when to_unsigned(83, 8) =>
			level <= to_unsigned(168, 8);
		when to_unsigned(84, 8) =>
			level <= to_unsigned(170, 8);
		when to_unsigned(85, 8) =>
			level <= to_unsigned(172, 8);
		when to_unsigned(86, 8) =>
			level <= to_unsigned(174, 8);
		when to_unsigned(87, 8) =>
			level <= to_unsigned(176, 8);
		when to_unsigned(88, 8) =>
			level <= to_unsigned(178, 8);
		when to_unsigned(89, 8) =>
			level <= to_unsigned(180, 8);
		when to_unsigned(90, 8) =>
			level <= to_unsigned(182, 8);
		when to_unsigned(91, 8) =>
			level <= to_unsigned(184, 8);
		when to_unsigned(92, 8) =>
			level <= to_unsigned(186, 8);
		when to_unsigned(93, 8) =>
			level <= to_unsigned(188, 8);
		when to_unsigned(94, 8) =>
			level <= to_unsigned(190, 8);
		when to_unsigned(95, 8) =>
			level <= to_unsigned(192, 8);
		when to_unsigned(96, 8) =>
			level <= to_unsigned(194, 8);
		when to_unsigned(97, 8) =>
			level <= to_unsigned(196, 8);
		when to_unsigned(98, 8) =>
			level <= to_unsigned(198, 8);
		when to_unsigned(99, 8) =>
			level <= to_unsigned(200, 8);
		when to_unsigned(100, 8) =>
			level <= to_unsigned(202, 8);
		when to_unsigned(101, 8) =>
			level <= to_unsigned(204, 8);
		when to_unsigned(102, 8) =>
			level <= to_unsigned(206, 8);
		when to_unsigned(103, 8) =>
			level <= to_unsigned(208, 8);
		when to_unsigned(104, 8) =>
			level <= to_unsigned(210, 8);
		when to_unsigned(105, 8) =>
			level <= to_unsigned(212, 8);
		when to_unsigned(106, 8) =>
			level <= to_unsigned(214, 8);
		when to_unsigned(107, 8) =>
			level <= to_unsigned(216, 8);
		when to_unsigned(108, 8) =>
			level <= to_unsigned(218, 8);
		when to_unsigned(109, 8) =>
			level <= to_unsigned(220, 8);
		when to_unsigned(110, 8) =>
			level <= to_unsigned(222, 8);
		when to_unsigned(111, 8) =>
			level <= to_unsigned(224, 8);
		when to_unsigned(112, 8) =>
			level <= to_unsigned(226, 8);
		when to_unsigned(113, 8) =>
			level <= to_unsigned(228, 8);
		when to_unsigned(114, 8) =>
			level <= to_unsigned(230, 8);
		when to_unsigned(115, 8) =>
			level <= to_unsigned(232, 8);
		when to_unsigned(116, 8) =>
			level <= to_unsigned(234, 8);
		when to_unsigned(117, 8) =>
			level <= to_unsigned(236, 8);
		when to_unsigned(118, 8) =>
			level <= to_unsigned(238, 8);
		when to_unsigned(119, 8) =>
			level <= to_unsigned(240, 8);
		when to_unsigned(120, 8) =>
			level <= to_unsigned(242, 8);
		when to_unsigned(121, 8) =>
			level <= to_unsigned(244, 8);
		when to_unsigned(122, 8) =>
			level <= to_unsigned(246, 8);
		when to_unsigned(123, 8) =>
			level <= to_unsigned(248, 8);
		when to_unsigned(124, 8) =>
			level <= to_unsigned(250, 8);
		when to_unsigned(125, 8) =>
			level <= to_unsigned(252, 8);
		when to_unsigned(126, 8) =>
			level <= to_unsigned(254, 8);
		when to_unsigned(127, 8) =>
			level <= to_unsigned(256, 8);
		when to_unsigned(128, 8) =>
			level <= to_unsigned(258, 8);
		when to_unsigned(129, 8) =>
			level <= to_unsigned(260, 8);
		when to_unsigned(130, 8) =>
			level <= to_unsigned(262, 8);
		when to_unsigned(131, 8) =>
			level <= to_unsigned(264, 8);
		when to_unsigned(132, 8) =>
			level <= to_unsigned(266, 8);
		when to_unsigned(133, 8) =>
			level <= to_unsigned(268, 8);
		when to_unsigned(134, 8) =>
			level <= to_unsigned(270, 8);
		when to_unsigned(135, 8) =>
			level <= to_unsigned(272, 8);
		when to_unsigned(136, 8) =>
			level <= to_unsigned(274, 8);
		when to_unsigned(137, 8) =>
			level <= to_unsigned(276, 8);
		when to_unsigned(138, 8) =>
			level <= to_unsigned(278, 8);
		when to_unsigned(139, 8) =>
			level <= to_unsigned(280, 8);
		when to_unsigned(140, 8) =>
			level <= to_unsigned(282, 8);
		when to_unsigned(141, 8) =>
			level <= to_unsigned(284, 8);
		when to_unsigned(142, 8) =>
			level <= to_unsigned(286, 8);
		when to_unsigned(143, 8) =>
			level <= to_unsigned(288, 8);
		when to_unsigned(144, 8) =>
			level <= to_unsigned(290, 8);
		when to_unsigned(145, 8) =>
			level <= to_unsigned(292, 8);
		when to_unsigned(146, 8) =>
			level <= to_unsigned(294, 8);
		when to_unsigned(147, 8) =>
			level <= to_unsigned(296, 8);
		when to_unsigned(148, 8) =>
			level <= to_unsigned(298, 8);
		when to_unsigned(149, 8) =>
			level <= to_unsigned(300, 8);
		when to_unsigned(150, 8) =>
			level <= to_unsigned(302, 8);
		when to_unsigned(151, 8) =>
			level <= to_unsigned(304, 8);
		when to_unsigned(152, 8) =>
			level <= to_unsigned(306, 8);
		when to_unsigned(153, 8) =>
			level <= to_unsigned(308, 8);
		when to_unsigned(154, 8) =>
			level <= to_unsigned(310, 8);
		when to_unsigned(155, 8) =>
			level <= to_unsigned(312, 8);
		when to_unsigned(156, 8) =>
			level <= to_unsigned(134, 8);
		when to_unsigned(157, 8) =>
			level <= to_unsigned(316, 8);
		when to_unsigned(158, 8) =>
			level <= to_unsigned(318, 8);
		when to_unsigned(159, 8) =>
			level <= to_unsigned(320, 8);
		when to_unsigned(160, 8) =>
			level <= to_unsigned(322, 8);
		when to_unsigned(161, 8) =>
			level <= to_unsigned(324, 8);
		when to_unsigned(162, 8) =>
			level <= to_unsigned(326, 8);
		when to_unsigned(163, 8) =>
			level <= to_unsigned(328, 8);
		when to_unsigned(164, 8) =>
			level <= to_unsigned(330, 8);
		when to_unsigned(165, 8) =>
			level <= to_unsigned(332, 8);
		when to_unsigned(166, 8) =>
			level <= to_unsigned(334, 8);
		when to_unsigned(167, 8) =>
			level <= to_unsigned(336, 8);
		when to_unsigned(168, 8) =>
			level <= to_unsigned(338, 8);
		when to_unsigned(169, 8) =>
			level <= to_unsigned(340, 8);
		when to_unsigned(170, 8) =>
			level <= to_unsigned(342, 8);
		when to_unsigned(171, 8) =>
			level <= to_unsigned(344, 8);
		when to_unsigned(172, 8) =>
			level <= to_unsigned(346, 8);
		when to_unsigned(173, 8) =>
			level <= to_unsigned(348, 8);
		when to_unsigned(174, 8) =>
			level <= to_unsigned(350, 8);
		when to_unsigned(175, 8) =>
			level <= to_unsigned(352, 8);
		when to_unsigned(176, 8) =>
			level <= to_unsigned(354, 8);
		when to_unsigned(177, 8) =>
			level <= to_unsigned(356, 8);
		when to_unsigned(178, 8) =>
			level <= to_unsigned(358, 8);
		when to_unsigned(179, 8) =>
			level <= to_unsigned(360, 8);
		when to_unsigned(180, 8) =>
			level <= to_unsigned(362, 8);
		when to_unsigned(181, 8) =>
			level <= to_unsigned(364, 8);
		when to_unsigned(182, 8) =>
			level <= to_unsigned(366, 8);
		when to_unsigned(183, 8) =>
			level <= to_unsigned(368, 8);
		when to_unsigned(184, 8) =>
			level <= to_unsigned(370, 8);
		when to_unsigned(185, 8) =>
			level <= to_unsigned(372, 8);
		when to_unsigned(186, 8) =>
			level <= to_unsigned(374, 8);
		when to_unsigned(187, 8) =>
			level <= to_unsigned(376, 8);
		when to_unsigned(188, 8) =>
			level <= to_unsigned(378, 8);
		when to_unsigned(189, 8) =>
			level <= to_unsigned(380, 8);
		when to_unsigned(190, 8) =>
			level <= to_unsigned(382, 8);
		when to_unsigned(191, 8) =>
			level <= to_unsigned(384, 8);
		when to_unsigned(192, 8) =>
			level <= to_unsigned(386, 8);
		when to_unsigned(193, 8) =>
			level <= to_unsigned(388, 8);
		when to_unsigned(194, 8) =>
			level <= to_unsigned(390, 8);
		when to_unsigned(195, 8) =>
			level <= to_unsigned(392, 8);
		when to_unsigned(196, 8) =>
			level <= to_unsigned(394, 8);
		when to_unsigned(197, 8) =>
			level <= to_unsigned(396, 8);
		when to_unsigned(198, 8) =>
			level <= to_unsigned(398, 8);
		when to_unsigned(199, 8) =>
			level <= to_unsigned(400, 8);
		when to_unsigned(200, 8) =>
			level <= to_unsigned(402, 8);
		when to_unsigned(201, 8) =>
			level <= to_unsigned(404, 8);
		when to_unsigned(202, 8) =>
			level <= to_unsigned(406, 8);
		when to_unsigned(203, 8) =>
			level <= to_unsigned(408, 8);
		when to_unsigned(204, 8) =>
			level <= to_unsigned(410, 8);
		when to_unsigned(205, 8) =>
			level <= to_unsigned(412, 8);
		when to_unsigned(206, 8) =>
			level <= to_unsigned(414, 8);
		when to_unsigned(207, 8) =>
			level <= to_unsigned(416, 8);
		when to_unsigned(208, 8) =>
			level <= to_unsigned(418, 8);
		when to_unsigned(209, 8) =>
			level <= to_unsigned(420, 8);
		when to_unsigned(210, 8) =>
			level <= to_unsigned(422, 8);
		when to_unsigned(211, 8) =>
			level <= to_unsigned(424, 8);
		when to_unsigned(212, 8) =>
			level <= to_unsigned(426, 8);
		when to_unsigned(213, 8) =>
			level <= to_unsigned(428, 8);
		when to_unsigned(214, 8) =>
			level <= to_unsigned(430, 8);
		when to_unsigned(215, 8) =>
			level <= to_unsigned(432, 8);
		when to_unsigned(216, 8) =>
			level <= to_unsigned(434, 8);
		when to_unsigned(217, 8) =>
			level <= to_unsigned(436, 8);
		when to_unsigned(218, 8) =>
			level <= to_unsigned(438, 8);
		when to_unsigned(219, 8) =>
			level <= to_unsigned(440, 8);
		when to_unsigned(220, 8) =>
			level <= to_unsigned(442, 8);
		when to_unsigned(221, 8) =>
			level <= to_unsigned(444, 8);
		when to_unsigned(222, 8) =>
			level <= to_unsigned(446, 8);
		when to_unsigned(223, 8) =>
			level <= to_unsigned(448, 8);
		when to_unsigned(224, 8) =>
			level <= to_unsigned(450, 8);
		when to_unsigned(225, 8) =>
			level <= to_unsigned(452, 8);
		when to_unsigned(226, 8) =>
			level <= to_unsigned(454, 8);
		when to_unsigned(227, 8) =>
			level <= to_unsigned(456, 8);
		when to_unsigned(228, 8) =>
			level <= to_unsigned(458, 8);
		when to_unsigned(229, 8) =>
			level <= to_unsigned(460, 8);
		when to_unsigned(230, 8) =>
			level <= to_unsigned(462, 8);
		when to_unsigned(231, 8) =>
			level <= to_unsigned(464, 8);
		when to_unsigned(232, 8) =>
			level <= to_unsigned(466, 8);
		when to_unsigned(233, 8) =>
			level <= to_unsigned(468, 8);
		when to_unsigned(234, 8) =>
			level <= to_unsigned(470, 8);
		when to_unsigned(235, 8) =>
			level <= to_unsigned(472, 8);
		when to_unsigned(236, 8) =>
			level <= to_unsigned(474, 8);
		when to_unsigned(237, 8) =>
			level <= to_unsigned(476, 8);
		when to_unsigned(238, 8) =>
			level <= to_unsigned(478, 8);
		
		when others =>
			level <= "00000000";
	end case;
end process;

end Behavioral;

